module pcalu (
    input wire [31:0] read1,
    output wire [31:0] out1,
    input wire CLK
);
endmodule
